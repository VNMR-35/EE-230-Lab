B6. RLC Bandpass Filter Vinamra Baghel 190010070
* <element-name> <nodes> <value/model>
l 1 2 10m
c 2 3 0.1u
r 3 0 1k
vin 1 0 dc 0 ac 1
*analysis command
.ac dec 10 1 10Meg
.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set xbrushwidth = 2
plot vdb(3) vdb(1)
meas ac peak MAX vmag(3)
meas ac fpeak WHEN vmag(3) = peak
let f3db = peak/sqrt(2)
meas ac f1 WHEN vmag(3)=f3db RISE=1
meas ac f2 WHEN vmag(3)=f3db FALL=1
.endc
.end
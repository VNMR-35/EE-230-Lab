Vinamra Baghel 190010070 Simulation of MOSFET Circuits

.model NXYAA5U nmos Level=1 Vto=0.7 KP=100u w=10u L=1u Gamma=0 Phi=0.65 Lambda=0.0

m d g 0 0 NXYAA5U
vg g 0 1.5
vd d 0 3

.op
.control
run
print -i(vd)
.endc
.end
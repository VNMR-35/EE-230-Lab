Vinamra Baghel 190010070 Common-Collector Amplifier: Midband Voltage Gain

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3 BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40 tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

*Netlist
rb c b 1M
re e gnd 10k
rs in in2 0
c1 in2 b 10u
c2 c out 10u
Q c b e bc547a
Vcc c gnd 12
Vin in gnd dc 0 ac sin()

*Analysis
.ac 

*Control
.control
run

.endc
.end
Vinamra Baghel 190010070 Full Wave Rectifier

.include ua741.txt
.include IN914.txt

*Netlist
r1 in neg1 10k
r2 neg1 in1 10k
rs1 in neg2 10k
rs2 in1 neg2 5k
rf neg2 out 10k
rl out gnd 1k
D1 o1 neg1 1N914
D2 in1 o1 1N914
X1 gnd neg1 pp np o1 ua741
X2 gnd neg2 pp np out ua741
Vccp pp gnd 12
Vccn np gnd -12
Vin in gnd sin(0 1 100 0 0 0)

*Analysis
.tran 1u 40m
.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set color4 = green
set xbrushwidth = 2
plot v(out) vs v(in)
.endc
.end
Vinamra Baghel 190010070 NMOS Current Mirror based Current Source

.model NXYAA5U nmos Level=1 Vto=1 KP=100u w=10u L=1u Gamma=0 Phi=0.65 Lambda=0.01

r dd g 8.2k
m1 g g 0 0 NXYAA5U
m2 o g 0 0 NXYAA5U
vo o 0 1
vdd dd 0 12

.dc vo 1 5 0.2
.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set color4 = green
set xbrushwidth = 2.5
*print i(vdd) i(vo)
plot i(vdd) i(vo)
.endc
.end
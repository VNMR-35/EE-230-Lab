Vinamra Baghel 190010070 Improved Half Wave Rectifier-A

.include ua741.txt
.include IN914.txt

*Netlist
r1 in neg 10k
r2 neg out 10k
rl out gnd 1k
D1 neg o1 1N914
D2 o1 out 1N914
X1 gnd neg pp np o1 ua741
Vccp pp gnd 12
Vccn np gnd -12
Vin in gnd sin(0 1 100 0 0 0)

*Analysis
.tran 1u 40m
.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set color4 = green
set xbrushwidth = 2
plot v(out) vs v(in)
.endc
.end
B1. RC Integrator Vinamra Baghel 190010070
* <element-name> <nodes> <value/model>
r 1 2 10k
c 2 0 0.1u
v 1 0 pulse(0 5 0.5m 0 0 10m 20m)
*analysis command
.tran 10u 100m
.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set xbrushwidth = 2
plot v(2) v(1)
.endc
.end
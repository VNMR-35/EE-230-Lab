B2. RC Differentiator Vinamra Baghel 190010070
* <element-name> <nodes> <value/model>
r 2 0 10k
c 1 2 0.1u
v 1 0 pulse(0 5 0 0 0 5m 10m)
*analysis command
.tran 10u 100m
.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set xbrushwidth = 2
plot v(2) v(1)
.endc
.end
Vinamra Baghel 190010070 Two Stage Amplifier: Biasing Circuit

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3 BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40 tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

*Netlist
rs in in2 0
r1 cc b1 10k
r2 b1 gnd 2.2k
rc cc c1 1.2k
re1 e1 gnd 1k
re2 de2 gnd 10k
rl out gnd 10k
cap1 in2 b1 10u
cape e1 gnd 100u
cap2 e2 out 10u
Q1 c1 b1 e1 bc547a
Q2 cc b2 e2 bc547a
vb2 c1 b2 0
ve2 e2 de2 0
Vcc cc gnd 12
Vin in gnd dc 0 ac 10m

*Analysis
.ac dec 10 10 10Meg

*Control
.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set xbrushwidth = 2
print v(out)*100
plot vdb(out)
.endc
.end
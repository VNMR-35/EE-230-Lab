Vinamra Baghel 190010070 Common-Collector Amplifier: Biasing Circuit

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3 BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40 tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

*Netlist
rb c db 1M
re de gnd 10k
Q c b e bc547a
ve e de 0
vb db b 0
Vcc c gnd 12

*Analysis
.op 

*Control
.control
run
print i(vb) i(ve) v(b) v(e)
.endc
.end
Vinamra Baghel 190010070 Wein Bridge Oscillator

.include ua741.txt

*Netlist
r1 gnd neg 4.7k
r2 neg out 10k
rs out 1 4.7k
cs 1 pos 0.1u
rp pos gnd 4.7k
cp pos gnd 0.1u
X1 pos neg pp np out ua741
Vccp pp gnd 12
Vccn np gnd -12

*Analysis
.tran 3u 270m 200m
.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set color4 = green
set xbrushwidth = 2
plot v(out)
.endc
.end
Vinamra Baghel 190010070 DC Power Supply with BJT Series Regulator

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3 BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40 tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f
.model SL100 NPN IS=100f BF=80 ISE=10.3f IKF=50m NE=1.3 BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=100 RE=1 RC=10 tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

.SUBCKT ZENER_12 1 2
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 10.8
.MODEL DF D (IS=27.5p RS=0.620 N=1.10 CJO=78.3p VJ=1.00 M=0.330 TT=50.1n)
.MODEL DR D (IS=5.49f RS=50 N=1.77)
.ENDS

*Netlist
Q1 in 1 out SL100
Q2 1 2 3 bc547a
X gnd 3 ZENER_12
rc in 1 1k
r1 out 2 14k
r2 2 gnd 11k
rl out gnd 1k
vin in gnd dc 20

*Analysis
.op

*Control
.control
run
print all
.endc
.end
Vinamra Baghel 190010070 Common-Emitter Amplifier: Biasing Circuit

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3 BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40 tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

*Netlist
r1 cc db 10k
r2 db gnd 2.2k
rc cc dc 1.2k
re e gnd 1k
Q c b e bc547a
vb db b 0
vc dc c 0
Vcc cc gnd 12

*Analysis
.op

*Control
.control
run
print i(vb) i(vc) v(b) v(c) v(e)
.endc
.end